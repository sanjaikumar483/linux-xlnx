module test(input a,b, output c);
nand NAND (c,a,b);
endmodule
